magic
tech sky130A
magscale 1 2
timestamp 1709819701
<< nwell >>
rect 320 992 330 1063
rect 268 694 330 992
rect 320 630 330 694
rect 255 568 330 630
rect 320 486 330 568
<< poly >>
rect 144 269 174 610
rect 268 250 298 630
<< metal1 >>
rect 92 906 138 996
rect 220 681 294 698
rect 226 660 294 681
rect 226 630 307 660
rect 226 182 268 250
rect 92 54 138 100
use grid  grid_0
timestamp 1709745296
transform 1 0 61 0 1 10
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_0
timestamp 1709745296
transform 1 0 159 0 1 175
box -73 -101 73 101
use sky130_fd_pr__pfet_01v8_52K3FE  sky130_fd_pr__pfet_01v8_52K3FE_0
timestamp 1709745296
transform 1 0 159 0 1 780
box -109 -212 109 212
use via_m1_p  via_m1_p_0
timestamp 1709818676
transform 1 0 255 0 1 182
box 6 0 64 68
use via_m1_p  via_m1_p_1
timestamp 1709818676
transform 1 0 262 0 1 630
box 6 0 64 68
<< labels >>
rlabel space 33 988 288 1031 1 vdd
rlabel metal1 34 6 289 49 1 vss
rlabel poly 144 250 174 630 1 in
rlabel space 268 234 298 648 1 out
<< end >>
