magic
tech sky130A
magscale 1 2
timestamp 1709783307
<< nwell >>
rect -334 485 -265 1062
rect 39 1060 91 1062
rect 54 485 91 1060
rect 411 947 414 1062
rect 411 485 414 523
rect -11 -559 672 -521
rect -4 -760 672 -559
rect -5 -983 673 -760
rect -11 -1034 673 -983
rect -11 -1098 672 -1034
<< nmos >>
rect 142 -284 172 -134
rect 498 -284 528 -134
<< pmos >>
rect 93 -972 123 -822
rect 189 -972 219 -822
rect 449 -972 479 -822
rect 545 -972 575 -822
<< ndiff >>
rect 84 -146 142 -134
rect 84 -272 96 -146
rect 130 -272 142 -146
rect 84 -284 142 -272
rect 172 -146 230 -134
rect 172 -272 184 -146
rect 218 -272 230 -146
rect 172 -284 230 -272
rect 440 -146 498 -134
rect 440 -272 452 -146
rect 486 -272 498 -146
rect 440 -284 498 -272
rect 528 -146 586 -134
rect 528 -272 540 -146
rect 574 -272 586 -146
rect 528 -284 586 -272
<< pdiff >>
rect 31 -834 93 -822
rect 31 -960 43 -834
rect 77 -960 93 -834
rect 31 -972 93 -960
rect 123 -834 189 -822
rect 123 -960 139 -834
rect 173 -960 189 -834
rect 123 -972 189 -960
rect 219 -834 281 -822
rect 219 -960 235 -834
rect 269 -960 281 -834
rect 219 -972 281 -960
rect 387 -834 449 -822
rect 387 -960 399 -834
rect 433 -960 449 -834
rect 387 -972 449 -960
rect 479 -834 545 -822
rect 479 -960 495 -834
rect 529 -960 545 -834
rect 479 -972 545 -960
rect 575 -834 637 -822
rect 575 -960 591 -834
rect 625 -960 637 -834
rect 575 -972 637 -960
<< ndiffc >>
rect 96 -272 130 -146
rect 184 -272 218 -146
rect 452 -272 486 -146
rect 540 -272 574 -146
<< pdiffc >>
rect 43 -960 77 -834
rect 139 -960 173 -834
rect 235 -960 269 -834
rect 399 -960 433 -834
rect 495 -960 529 -834
rect 591 -960 625 -834
<< psubdiff >>
rect 33 -79 57 -45
rect 257 -79 281 -45
rect 389 -79 413 -45
rect 613 -79 637 -45
<< nsubdiff >>
rect 32 -1027 280 -1026
rect 32 -1061 81 -1027
rect 228 -1061 280 -1027
rect 32 -1062 280 -1061
rect 388 -1027 636 -1026
rect 388 -1061 437 -1027
rect 584 -1061 636 -1027
rect 388 -1062 636 -1061
<< psubdiffcont >>
rect 57 -79 257 -45
rect 413 -79 613 -45
<< nsubdiffcont >>
rect 81 -1061 228 -1027
rect 437 -1061 584 -1027
<< poly >>
rect 142 -134 172 -108
rect 498 -134 528 -108
rect 2 -297 60 -279
rect 2 -331 14 -297
rect 48 -331 60 -297
rect 142 -322 172 -284
rect 254 -298 312 -280
rect 2 -347 60 -331
rect 129 -340 187 -322
rect 15 -678 64 -347
rect 129 -374 141 -340
rect 175 -374 187 -340
rect 254 -332 266 -298
rect 300 -332 312 -298
rect 254 -348 312 -332
rect 358 -297 416 -279
rect 358 -331 370 -297
rect 404 -331 416 -297
rect 498 -322 528 -284
rect 610 -298 668 -280
rect 358 -347 416 -331
rect 485 -340 543 -322
rect 129 -390 187 -374
rect 2 -696 60 -678
rect 2 -730 14 -696
rect 48 -730 60 -696
rect 2 -746 60 -730
rect 127 -684 185 -666
rect 248 -678 300 -348
rect 371 -678 420 -347
rect 485 -374 497 -340
rect 531 -374 543 -340
rect 610 -332 622 -298
rect 656 -332 668 -298
rect 610 -348 668 -332
rect 485 -390 543 -374
rect 248 -679 312 -678
rect 127 -718 139 -684
rect 173 -718 185 -684
rect 127 -734 185 -718
rect 254 -696 312 -679
rect 254 -730 266 -696
rect 300 -730 312 -696
rect 142 -777 172 -734
rect 254 -746 312 -730
rect 358 -696 416 -678
rect 358 -730 370 -696
rect 404 -730 416 -696
rect 358 -746 416 -730
rect 483 -684 541 -666
rect 604 -678 656 -348
rect 604 -679 668 -678
rect 483 -718 495 -684
rect 529 -718 541 -684
rect 483 -734 541 -718
rect 610 -696 668 -679
rect 610 -730 622 -696
rect 656 -730 668 -696
rect 498 -777 528 -734
rect 610 -746 668 -730
rect 93 -807 219 -777
rect 93 -822 123 -807
rect 189 -822 219 -807
rect 449 -807 575 -777
rect 449 -822 479 -807
rect 545 -822 575 -807
rect 93 -998 123 -972
rect 189 -998 219 -972
rect 449 -998 479 -972
rect 545 -998 575 -972
<< polycont >>
rect 14 -331 48 -297
rect 141 -374 175 -340
rect 266 -332 300 -298
rect 370 -331 404 -297
rect 14 -730 48 -696
rect 497 -374 531 -340
rect 622 -332 656 -298
rect 139 -718 173 -684
rect 266 -730 300 -696
rect 370 -730 404 -696
rect 495 -718 529 -684
rect 622 -730 656 -696
<< locali >>
rect 96 -146 130 -130
rect 2 -297 60 -279
rect 96 -288 130 -272
rect 184 -146 218 -130
rect 184 -288 218 -272
rect 452 -146 486 -130
rect 2 -331 14 -297
rect 48 -331 60 -297
rect 254 -298 312 -280
rect 2 -347 60 -331
rect 129 -340 187 -322
rect 129 -374 141 -340
rect 175 -374 187 -340
rect 254 -332 266 -298
rect 300 -332 312 -298
rect 254 -348 312 -332
rect 358 -297 416 -279
rect 452 -288 486 -272
rect 540 -146 574 -130
rect 540 -288 574 -272
rect 358 -331 370 -297
rect 404 -331 416 -297
rect 610 -298 668 -280
rect 358 -347 416 -331
rect 485 -340 543 -322
rect 129 -390 187 -374
rect 485 -374 497 -340
rect 531 -374 543 -340
rect 610 -332 622 -298
rect 656 -332 668 -298
rect 610 -348 668 -332
rect 485 -390 543 -374
rect 2 -696 60 -678
rect 2 -730 14 -696
rect 48 -730 60 -696
rect 2 -746 60 -730
rect 127 -684 185 -666
rect 127 -718 139 -684
rect 173 -718 185 -684
rect 127 -734 185 -718
rect 254 -696 312 -678
rect 254 -730 266 -696
rect 300 -730 312 -696
rect 254 -746 312 -730
rect 358 -696 416 -678
rect 358 -730 370 -696
rect 404 -730 416 -696
rect 358 -746 416 -730
rect 483 -684 541 -666
rect 483 -718 495 -684
rect 529 -718 541 -684
rect 483 -734 541 -718
rect 610 -696 668 -678
rect 610 -730 622 -696
rect 656 -730 668 -696
rect 610 -746 668 -730
rect 43 -834 77 -818
rect 43 -976 77 -960
rect 139 -834 173 -818
rect 139 -976 173 -960
rect 235 -834 269 -818
rect 235 -976 269 -960
rect 399 -834 433 -818
rect 399 -976 433 -960
rect 495 -834 529 -818
rect 495 -976 529 -960
rect 591 -834 625 -818
rect 591 -976 625 -960
rect 23 -1023 289 -1019
rect 23 -1066 29 -1023
rect 284 -1066 289 -1023
rect 23 -1069 289 -1066
rect 379 -1023 645 -1019
rect 379 -1066 385 -1023
rect 640 -1066 645 -1023
rect 379 -1069 645 -1066
<< viali >>
rect 30 -45 285 -41
rect 30 -79 57 -45
rect 57 -79 257 -45
rect 257 -79 285 -45
rect 30 -84 285 -79
rect 386 -45 641 -41
rect 386 -79 413 -45
rect 413 -79 613 -45
rect 613 -79 641 -45
rect 386 -84 641 -79
rect 96 -272 130 -146
rect 184 -272 218 -146
rect 452 -272 486 -146
rect 14 -331 48 -297
rect 141 -374 175 -340
rect 266 -332 300 -298
rect 540 -272 574 -146
rect 370 -331 404 -297
rect 497 -374 531 -340
rect 622 -332 656 -298
rect 14 -730 48 -696
rect 139 -718 173 -684
rect 266 -730 300 -696
rect 370 -730 404 -696
rect 495 -718 529 -684
rect 622 -730 656 -696
rect 43 -960 77 -834
rect 139 -960 173 -834
rect 235 -960 269 -834
rect 399 -960 433 -834
rect 495 -960 529 -834
rect 591 -960 625 -834
rect 29 -1027 284 -1023
rect 29 -1061 81 -1027
rect 81 -1061 228 -1027
rect 228 -1061 284 -1027
rect 29 -1066 284 -1061
rect 385 -1027 640 -1023
rect 385 -1061 437 -1027
rect 437 -1061 584 -1027
rect 584 -1061 640 -1027
rect 385 -1066 640 -1061
<< metal1 >>
rect 18 -41 297 -35
rect 18 -84 30 -41
rect 285 -84 297 -41
rect 18 -90 297 -84
rect 374 -41 653 -35
rect 374 -84 386 -41
rect 641 -84 653 -41
rect 374 -90 653 -84
rect 90 -146 136 -134
rect 90 -238 96 -146
rect 2 -272 96 -238
rect 130 -272 136 -146
rect 2 -284 136 -272
rect 178 -146 224 -134
rect 178 -272 184 -146
rect 218 -238 224 -146
rect 446 -146 492 -134
rect 446 -238 452 -146
rect 218 -272 312 -238
rect 178 -284 312 -272
rect 2 -297 60 -284
rect 2 -331 14 -297
rect 48 -331 60 -297
rect 254 -298 312 -284
rect 2 -347 60 -331
rect 129 -340 187 -322
rect 129 -374 141 -340
rect 175 -374 187 -340
rect 254 -332 266 -298
rect 300 -332 312 -298
rect 254 -348 312 -332
rect 358 -272 452 -238
rect 486 -272 492 -146
rect 358 -284 492 -272
rect 534 -146 580 -134
rect 534 -272 540 -146
rect 574 -238 580 -146
rect 574 -272 668 -238
rect 534 -284 668 -272
rect 358 -297 416 -284
rect 358 -331 370 -297
rect 404 -331 416 -297
rect 610 -298 668 -284
rect 358 -347 416 -331
rect 485 -340 543 -322
rect 129 -390 187 -374
rect 485 -374 497 -340
rect 531 -374 543 -340
rect 610 -332 622 -298
rect 656 -332 668 -298
rect 610 -348 668 -332
rect 485 -390 543 -374
rect 2 -696 60 -678
rect 2 -730 14 -696
rect 48 -730 60 -696
rect 2 -822 60 -730
rect 127 -684 185 -666
rect 127 -718 139 -684
rect 173 -718 185 -684
rect 127 -734 185 -718
rect 254 -696 312 -678
rect 254 -730 266 -696
rect 300 -730 312 -696
rect 254 -822 312 -730
rect 2 -834 83 -822
rect 2 -863 43 -834
rect 37 -960 43 -863
rect 77 -960 83 -834
rect 37 -972 83 -960
rect 133 -834 179 -822
rect 133 -960 139 -834
rect 173 -960 179 -834
rect 133 -972 179 -960
rect 229 -834 312 -822
rect 229 -960 235 -834
rect 269 -880 312 -834
rect 358 -696 416 -678
rect 358 -730 370 -696
rect 404 -730 416 -696
rect 358 -822 416 -730
rect 483 -684 541 -666
rect 483 -718 495 -684
rect 529 -718 541 -684
rect 483 -734 541 -718
rect 610 -696 668 -678
rect 610 -730 622 -696
rect 656 -730 668 -696
rect 610 -822 668 -730
rect 358 -834 439 -822
rect 358 -863 399 -834
rect 269 -960 275 -880
rect 229 -972 275 -960
rect 393 -960 399 -863
rect 433 -960 439 -834
rect 393 -972 439 -960
rect 489 -834 535 -822
rect 489 -960 495 -834
rect 529 -960 535 -834
rect 489 -972 535 -960
rect 585 -834 668 -822
rect 585 -960 591 -834
rect 625 -880 668 -834
rect 625 -960 631 -880
rect 585 -972 631 -960
rect 17 -1023 296 -1017
rect 17 -1066 29 -1023
rect 284 -1066 296 -1023
rect 17 -1072 296 -1066
rect 373 -1023 652 -1017
rect 373 -1066 385 -1023
rect 640 -1066 652 -1023
rect 373 -1072 652 -1066
use inverter_ahorasi  inverter_ahorasi_0
timestamp 1709782608
transform 1 0 660 0 -1 -38
box 0 0 330 1063
use inverter_ahorasi  inverter_ahorasi_1
timestamp 1709782608
transform 1 0 -654 0 1 -1
box 0 0 330 1063
use nor  nor_0
timestamp 1709782608
transform -1 0 -11 0 -1 -35
box -7 0 639 1063
use nor  nor_1
timestamp 1709782608
transform 1 0 414 0 1 -1
box -7 0 639 1063
use pass_gate  pass_gate_0
timestamp 1709782608
transform 1 0 -265 0 1 -1
box -1 0 321 1063
use pass_gate  pass_gate_1
timestamp 1709782608
transform 1 0 91 0 1 -1
box -1 0 321 1063
<< labels >>
rlabel metal1 17 -1072 296 -1017 5 VDD
rlabel metal1 373 -1072 652 -1017 5 VDD
rlabel metal1 374 -90 653 -35 5 VSS
rlabel metal1 18 -90 297 -35 5 VSS
<< end >>
