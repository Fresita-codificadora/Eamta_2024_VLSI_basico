magic
tech sky130A
timestamp 1709780221
<< poly >>
rect 3 26 32 34
rect 3 9 9 26
rect 26 9 32 26
rect 3 0 32 9
<< polycont >>
rect 9 9 26 26
<< locali >>
rect 3 26 32 34
rect 3 9 9 26
rect 26 9 32 26
rect 3 0 32 9
<< viali >>
rect 9 9 26 26
<< metal1 >>
rect 3 26 32 34
rect 3 9 9 26
rect 26 9 32 26
rect 3 0 32 9
<< end >>
